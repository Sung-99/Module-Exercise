module ANDDd (
    input  A,     // First input
    input  B,     // Second input
    output  Y     // Output
);

	
	
	assign Y = A & B; // AND operation
	

endmodule